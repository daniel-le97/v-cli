module utils

struct Logger {
	name  string
	level string
}
